module datapath_tb;
    $display("test passed");
endmodule